module hammingEncoder_tb;
	reg [3:0] message;
	wire [6:0] codeword;
	
	hammingEncoder uut(.message(message), .codeword(codeword));
	
	initial begin
		message = 4'b0000; #10;
		message = 4'b0001; #10;
		message = 4'b0010; #10;
		message = 4'b0011; #10;
		message = 4'b0100; #10;
		message = 4'b0101; #10;
		message = 4'b0110; #10;
		message = 4'b0111; #10;
		message = 4'b1000; #10;
		message = 4'b1001; #10;
		message = 4'b1010; #10;
		message = 4'b1011; #10;
		message = 4'b1100; #10;
		message = 4'b1101; #10;
		message = 4'b1110; #10;
		message = 4'b1111; #10;
		$stop;
	end
	initial
		$monitor($time,": message = %b, codeword = %b",message, codeword);
endmodule